module Display( );



endmodule
