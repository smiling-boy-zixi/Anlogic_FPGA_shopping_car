module my_rxd( );



endmodule
