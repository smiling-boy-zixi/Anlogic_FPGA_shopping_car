`timescale 1ns/1ns

// Define colors RGB--8|8|8
`define RED		24'hFF0000 
`define GREEN	24'h00FF00 
`define BLUE  	24'h0000FF 
`define WHITE 	24'hFFFFFF 
`define BLACK 	24'h000000 
`define YELLOW	24'hFFFF00 
`define CYAN  	24'hFF00FF 
`define ROYAL 	24'h00FFFF 


module Display_2
#(
	parameter H_DISP = 640, //Resolution
	parameter V_DISP = 480

)
( 
	input  wire	 		clk,	
	input  wire			rst_n,	
	input  wire	[11:0]	lcd_xpos,	//lcd horizontal coordinate
	input  wire	[11:0]	lcd_ypos,	//lcd vertical coordinate
	
	output reg  [23:0]	lcd_data	//lcd data
);

//************************************
	parameter POS_X = 240;   //�ַ�������ʼ�������
	parameter POS_Y = 174;	 //�ַ�������ʼ��������
	parameter WIDTH = 160;
	parameter HEIGHT = 68;
	reg  [159:0] char[68:0]; 
	wire [11:0] x_cnt;    //counter
	wire [11:0] y_cnt;
	assign x_cnt = lcd_xpos - POS_X; //���ص�������ַ�������ʼ��ˮƽ����
	assign y_cnt = lcd_ypos - POS_Y; //���ص�������ַ�������ʼ����ֱ����
////**************************************
//	parameter POS_X_1 = 284;		//�ڶ��������ַ�
//	parameter POS_Y_1 = 256;
//	parameter WIDTH_1   = 128;
//	parameter HEIGHT_1  = 32;
//	reg  [127:0] char_1[31:0];
//	wire [11:0] x_cnt_1;
//	wire [11:0] y_cnt_1;
//	assign x_cnt_1 = lcd_xpos - POS_X_1;
//	assign y_cnt_1 = lcd_xpos - POS_Y_1;

`ifdef VGA_TuDou
always@(posedge clk)
begin
	char[0]  <= 160'h0000000000000000000000000000000000000000;
	char[1]  <= 160'h0000000000000000000000000000000000000000;
	char[2]  <= 160'h0003800000000000000000000000000000000000;
	char[3]  <= 160'h0003C00000000060000000000000000000000080;
	char[4]  <= 160'h0003C0000FFFFFF0000000000000000003FFFFC0;
	char[5]  <= 160'h0003C00000000000000000000000000000000000;
	char[6]  <= 160'h0003C0000000000000000000000007E000000000;
	char[7]  <= 160'h0003C00000000000000000000000083800000000;
	char[8]  <= 160'h0003C00000000000000000000000101800000000;
	char[9]  <= 160'h0003C00001000080000000000000200C00000000;	
	char[10] <= 160'h0003C00001FFFFC0000000000000200C00000000;
	char[11] <= 160'h07FFC3800300C000000000000000018000000030;
	char[12] <= 160'h0003C0F001800180000000000000300C1FFFFFF8;
	char[13] <= 160'h1FFFFFF801800180000000000000000C000C3000;
	char[14] <= 160'h0C03C00001800180000000000000001800083000;
	char[15] <= 160'h0003C00001800180000000000000001800183000;
	char[16] <= 160'h0003C00001800180000000000000003000183000;
	char[17] <= 160'h0003C00001FFFF80000000000000006000183000;
	char[18] <= 160'h0003C0000180018000000000000000C000183000;
	char[19] <= 160'h0003C00001000000000000000000018000183000;
	char[20] <= 160'h0003C00000400400000000000000030000303008;
	char[21] <= 160'h0003C00000200F00000000000000020000303008;
	char[22] <= 160'h0003C00000300E00000000000000040400303008;
	char[23] <= 160'h0003C00000180C00000000000000080400603008;
	char[24] <= 160'h0003C00000181800000000000000100400603008;
	char[25] <= 160'h0003C01800181000000000000000200C00C03008;	
	char[26] <= 160'h0003C03C001830000000000000003FF80180301C;
	char[27] <= 160'h7FFFFFFE000020180000000000003FF803003FFC;
	char[28] <= 160'h300000003FFFFFFC000000000000000006001FF8;
	char[29] <= 160'h0000000000000000000000000000000018000000;
	char[30] <= 160'h0000000000000000000000000000000020000000;
	char[31] <= 160'h0000000000000000000000000000000000000000;
	//*********************************************************	
	char[32] <= 160'h0000000000000000000000000000000000000000;
	char[33] <= 160'h0000000000000000000000000000000000000000;
	char[34] <= 160'h0000000000000000000000000000000000000000;
	char[35] <= 160'h0000000000000000000000000000000000000000;
	//*******************************************************
	char[36] <= 160'h0000000000000000000000000000000000000000;//1
	char[37] <= 160'h0000000000000000000000000000000000000000;//2
	char[38] <= 160'h000000402000000100000080000000000C000000;//3
	char[39] <= 160'h0000006038000001800000E4004001000E000000;//4
	char[40] <= 160'h0000004030000001800000C7FFE003800C100000;//5
	char[41] <= 160'h0000004030000001818001C6004003030C180000;//6
	char[42] <= 160'h00000040300007FFFFC00186004003018C300000;//7
	char[43] <= 160'h0000004C308000018000018600400618CC200000;//8
	char[44] <= 160'h00001FFEFFC0000180000306004007FCCC400000;//9
	char[45] <= 160'h00000041308000018010030600400400CCC00000;//10	
	char[46] <= 160'h0000004031801FFFFFF8020600400C004C800000;//11
	char[47] <= 160'h000000403180000000380706004008020C100000;//12
	char[48] <= 160'h000000463180004040200707FFC00811FFF80000;//13
	char[49] <= 160'h000000792180003070400F0618401FF900300000;//14
	char[50] <= 160'h000001C0E180001860000B001800130100300000;//15
	char[51] <= 160'h00001F4061800018600013001800230100300000;//16
	char[52] <= 160'h00003840788804086000330018000301FFF00000;//17
	char[53] <= 160'h00001040DCC80308600023061800031900300000;//18
	char[54] <= 160'h000000408CC801804000030618303FF900300000;//19
	char[55] <= 160'h00000041046800C0400003041FF8030100300000;//20
	char[56] <= 160'h000007C2047800C0C01003041800030100300000;//21
	char[57] <= 160'h000001C4003C0080C038030C18000301FFF00000;//22
	char[58] <= 160'h00000088000C7FFFFFFC030C1800030100300000;//23
	char[59] <= 160'h00000200008000008000030E1800030100300000;//24
	char[60] <= 160'h0000021020400001C00003091800031100300000;//25
	char[61] <= 160'h0000060830600003380003199800036100300000;//26
	char[62] <= 160'h0000040C1830000607000310780003C100300000;//27
	char[63] <= 160'h00000C0C1830001801E003303800038100300000;//28
	char[64] <= 160'h00001C0C18300070007003200FFC030101F00000;//29
	char[65] <= 160'h00001808101003800030034001F8010100700000;//30
	char[66] <= 160'h0000000000003C00001002800000000100400000;//31
	char[67] <= 160'h0000000000000000000000000000000000000000;//32		
end

always@(posedge clk or negedge rst_n)//one
begin
	if(!rst_n)
		lcd_data <= 24'h0;
	else
	begin
		if((lcd_xpos >= POS_X) && (lcd_xpos  < POS_X + WIDTH)&&
		(lcd_ypos >= POS_Y)&&(lcd_ypos < POS_Y + HEIGHT))
		begin
			if(char[y_cnt][159 - x_cnt])
				lcd_data <= `BLACK;
			else
				lcd_data <= `WHITE;
		end
		else
			lcd_data <= `WHITE;
	end
end
`endif

endmodule